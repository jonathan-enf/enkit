module sub0;
  `include "common.svh"
endmodule : sub0
